library verilog;
use verilog.vl_types.all;
entity \MAC_\ is
    port(
        a               : in     vl_logic_vector(3 downto 0);
        b               : in     vl_logic_vector(3 downto 0);
        c               : in     vl_logic_vector(11 downto 0);
        result          : out    vl_logic_vector(11 downto 0);
        cout            : out    vl_logic
    );
end \MAC_\;
