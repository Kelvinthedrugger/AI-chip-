`include "MAC_4bit.v"
`include "HA.v"
`include "FA.v"
module MAC_8bit (
    input   [7:0]   a,
    input   [7:0]   b,
    input   [23:0]  c,
    output  [23:0]  result,
    output          cout
);

/* Here is your code */

endmodule




